b0VIM 8.2      �[]`    �  hermo                                   DESKTOP-BG953FA                         C:/Users/hermo/Develop/ped/pedropp/bet/app.py                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                utf-8 3210#"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     tp �      x            H   y                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              ad          x   �  �  �  �  �  �  �  �  (        �  �  �  �  ?  >  *    �  �  �  �  �  �  �  �  �  �  v  k  A  @  ?  >      �  �  �  �  y  x  `  ?  #    �  �  �  �  i  X  3    �
  ~
  R
  
  �	  �	  �	  Z	  .	  �  �  �  o  P      �  �  �  �  �  �  �  k  C    �  �  �  b  T  %    �  �  �  y  A    �  �  �  z  y  x  w  =  -    �  �  �  c  A       �  �  �  �  �  N                              def rec(user): @app.route('/recargas', methods=['GET', 'POST']) @app.route('/recargas/<user>', methods=['GET', 'POST'])               return render_template('fail.html', error = fallas['nolog'])         else:             return render_template('dashboard.html', user=user)              #flash('Bienvenido')             #enrutado a dashboard         if session['auth'] == 1 and session['name'] == user:     else:         return render_template('fail.html', error=fallas['noacces'])     if user == plantilla[0][1]:     plantilla = bd.leertodo() def dash(user): @app.route('/dashboard/<user>',  methods=['GET', 'POST'])            return render_template('registro.html')     else:                 return render_template('registro.html')                 flash("Datos ya existen")             except sqlite3.IntegrityError:                 return render_template('registro.html')             except ValueError:                 return redirect(url_for('log'))                 flash("registro realizado")                 bd.crear(datos)             try:             datos = (nombre, correo, password)         else:             return render_template('registro.html')             flash("No hay datos")         if nombre =="" or correo=="" or password =="":         password = request.form['password']         correo = request.form['correo']         nombre = request.form['nombre']     if request.method == 'POST':     #enrutado a registro def reg(): @app.route('/registro', methods=['GET', 'POST'])            return render_template('login.html')     else:                 return render_template('login.html')             except ValueError:                     return redirect(url_for('log'))                     flash("Datos Incorrectos")                 else:                         return redirect(url_for('dash', user=nombre))                         flash('Bienvenido')                         bd.log(str(nombre))                         #flash("te haz logeado correctamente")                         session['auth'] = 1                     else:                         return redirect(url_for('layad', user=nombre))                         flash('Bienvenido')                         session['auth'] = 1                     if nombre== str(plantilla[0][1]) and password == str(plantilla[0][3]):                     plantilla = bd.leertodo()                 if bd.existe(datos):             try:             datos = (nombre, password)         else:             return render_template('login.html')             flash("No hay datos")         if nombre =="" or password =="":                  session['auth'] = 0         session['name'] = nombre         session.clear()          password = request.form['password']         nombre = request.form['nombre']     if request.method == 'POST':      #enrutado a login def log(): @app.route('/login', methods=['GET', 'POST'])        return render_template('layout.html') def lay(): @app.route('/layout')        return render_template('index.html')     #enrutado a pagina inicial def hello(): @app.route('/')       session.permanent = True def session_manager(): @app.before_request  fallas = {'nolog':'Usuario no esta Logueado', 'noacces':'Usuario sin acceso a esta area'}  app.config.update(SESSION_COOKIE_SAMESITE="lax") app.secret_key="secretoenlamontana" app = Flask(__name__)  import bd import flask_wtf as wtf from flask import Flask, escape, request, render_template, url_for, redirect, flash, session, jsonify    #fecha 07/01/2021 11:07 PM # GP System C.A. #Author Luis Hermoso # _*_ coding: utf-8 _*_ #! usr\bin\env python ad  V  �	     H   �  �  �  >  =  <  ;    �  �  �  �  �  �  {  a  C  #  �  �  �  e  d  �  �  �  �  �  �  �  �  e  F  2    �  �  �  �  �  �  �  �  �  ^  ]  \  [  Z  /  #  �
  �
  �
  �
  �
  l
  R
  Q
  P
  O
  N
  9
  ,
  
  �	  �	  �	  �	  �	  �	  �	  w	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     app.run(host='     app.run(host='0.0.0.0', debug=1) if __name__ == '__main__':         return render_template('lista.html', plantilla = plantilla)     plantilla = bd.leertodo() def lista(): @app.route('/lista')         return jsonify(datos)             datos = bd.counteo()     elif datos == 'cuenta':         return jsonify(datos)         datos = bd.leertodo()     if datos == 'todo':     datos = request.args.get('datos') def json(): @app.route('/api/datos/', methods=['GET'])         return render_template('fail.html', error=fail) def fail(fail): @app.route('/fail')         return redirect(url_for('hello'))     cuenta = bd.counteo()     session['auth'] = 0     session['name'] = 'unknown'     session.clear()     bd.logout(session['name'])     #print(session['name']) def logout(): @app.route('/logout')                return render_template('fail.html', error=fallas['noacces'])         else:             return render_template('dashboard1.html', user=user, plantilla=plantilla, cuenta=cuenta)              #flash('Bienvvenido')         if session['auth'] == 1 and session['name'] == str(plantilla[0][1]):     else:         return render_template('fail.html', error=fallas['noacces'])     if user != plantilla[0][1]:     plantilla = bd.leertodo()     cuenta = bd.counteo() def layad(user): @app.route('/dashboard1/<user>', methods=['GET', 'POST'])        return render_template('documentacion.html') def doc(): @app.route('/documentacion', methods=['GET', 'POST'])            return render_template('fail.html', error=fallas['nolog'])     else:         return render_template('recargas.html', user=user)     if session['auth'] == 1 and  session['name'] == user: 